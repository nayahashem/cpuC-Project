`define W 4
`define PC 0

`define prog_size 8
`define Nplus 7
`define Nminus 2
`define Nmul 4
`define Nles 1
`define Nop `Nplus + `Nminus + `Nmul + `Nles

`define Nreg 3
`define Nconst 7
`define Nmem 1
`define Nmux 1

`define M 256 // memory size

`define CONST_FILE ",my_const.mem"
`define PROGRAM_FILE "my_program.mem"
