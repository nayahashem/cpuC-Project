`define W 4
`define PC 0

`define prog_size 8
`define Nplus 7
`define Nminus 6
`define Nmul 6
`define Nles 1
`define Nequ 6
`define Nop `Nplus + `Nminus + `Nmul + `Nles + `Nequ

`define Nreg 23
`define Nconst 24
`define Nmem 1
`define Nmux 6

`define M 256 // memory size

`define CONST_FILE ",my_const.mem"
`define PROGRAM_FILE "my_program.mem"
